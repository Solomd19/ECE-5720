`timescale 1ns/1ns

module tb_sixteen_bit_carry_lookahead_adder();

	//Inputs
	logic [15:0] X;
	logic [15:0] Y;
	logic Ci;
	
	//Outputs
	logic [15:0] S;
	logic Co;

	sixteen_bit_carry_lookahead_adder UUT(X, Y, Ci, S, Co);	

	initial
		begin
			X <= 16'b0000_0000_0000_0000;
			Y <= 16'b0000_0000_0000_0000;
			Ci <= 0;
			#10
			X <= 16'b0000_0000_0000_0001;
			Y <= 16'b0000_0000_0000_0000;
			#10
			X <= 16'b0000_0000_0000_0000;
			Y <= 16'b0000_0000_0000_0001;
			#10
			X <= 16'b0000_0000_0000_0001;
			Y <= 16'b0000_0000_0000_0001;
			#10
			X <= 16'b0000_0000_0000_0001;
			Y <= 16'b0000_0000_0000_0000;
			Ci <= 1;
			#10
			X <= 16'b0000_0000_0000_0000;
			Y <= 16'b0000_0000_0000_0001;
			#10
			X <= 16'b0000_0000_0000_0001;
			Y <= 16'b0000_0000_0000_0001;
			#10
			X <= 16'b1000_0000_0000_0000;
			Y <= 16'b0000_0000_0000_0000;
			#10
			X <= 16'b0000_0000_0000_0000;
			Y <= 16'b1000_0000_0000_0000;
			#10
			X <= 16'b1000_0000_0000_0000;
			Y <= 16'b1000_0000_0000_0000;
			#10
			X <= 16'b0000_0000_0000_0010;
			Y <= 16'b0000_0000_0000_0010;
			#10
			X <= 16'b0000_0000_0000_0100;
			Y <= 16'b0000_0000_0000_0100;
			#10
			X <= 16'b0000_0000_0000_1000;
			Y <= 16'b0000_0000_0000_1000;
			#10
			X <= 16'b1111_1111_1111_1111;
			Y <= 16'b1111_1111_1111_1111;
			Ci <= 1;
			#10
			$stop;
		end
endmodule
